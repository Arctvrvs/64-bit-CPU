// riscv_soc_4core.sv - Top level SoC placeholder

// Parameters: none
// Inputs: see port list below
// Outputs: see port list below

(* clock_gating_cell = "yes" *)
module riscv_soc_4core (
    input logic clk,
    input logic rst_n
);

    // Four core tiles and mesh would be instantiated here

endmodule
