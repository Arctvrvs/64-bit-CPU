// vector_fma512.sv - 512-bit vector fused multiply-add unit
//
// Purpose: Executes vector FMA operations across eight 64-bit lanes.
// Placeholder 5-stage pipeline producing results after five cycles.

// Parameters: none
// Inputs: see port list below
// Outputs: see port list below

(* clock_gating_cell = "yes" *)
module vector_fma512 (
    input  logic        clk,
    input  logic        rst_n,
    input  logic        valid_i,
    input  logic [511:0] src1_i,
    input  logic [511:0] src2_i,
    input  logic [511:0] src3_i,
    input  logic [63:0]  mask_i,
    output logic        valid_o,
    output logic [511:0] result_o
);

    localparam int STAGES = 5;
    logic [STAGES-1:0]        val_pipe;
    logic [511:0]             res_pipe [STAGES-1:0];

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            val_pipe <= '0;
        end else begin
            val_pipe[0] <= valid_i;
            for (int lane = 0; lane < 8; lane++) begin
                logic [63:0] a = src1_i[lane*64 +: 64];
                logic [63:0] b = src2_i[lane*64 +: 64];
                logic [63:0] c = src3_i[lane*64 +: 64];
                logic [63:0] prod = a * b + c;
                if (mask_i[lane])
                    res_pipe[0][lane*64 +: 64] <= prod;
                else
                    res_pipe[0][lane*64 +: 64] <= c;
            end
            for (int i = 1; i < STAGES; i++) begin
                val_pipe[i] <= val_pipe[i-1];
                res_pipe[i] <= res_pipe[i-1];
            end
        end
    end

    assign valid_o  = val_pipe[STAGES-1];
    assign result_o = res_pipe[STAGES-1];

endmodule
