// core_tile_2smts_8wide.sv - Placeholder dual-SMT core tile

// Parameters: none
// Inputs: see port list below
// Outputs: see port list below

(* clock_gating_cell = "yes" *)
module core_tile_2smts_8wide (
    input logic clk,
    input logic rst_n
);

    // submodules would be instantiated here in the future

endmodule
